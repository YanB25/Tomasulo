`timescale 1ns/1ps
`include "head.v"

module StoreStation(
    input clk,
    input 
)